`timescale 1ns / 1ps

module bin_count #(parameter MAX_COUNT = 255, WIDTH = 8)
(
	input rst, clk, cen,
	output [WIDTH-1:0] val
);
	//module description here
endmodule
